module uart
(
	
);


endmodule