module uart
(
	
);

endmodule
