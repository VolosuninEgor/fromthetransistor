module uart
(
	
);

endmodule